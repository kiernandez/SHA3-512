module tbkeccakP;

/////////////////////////////////////////

parameter inClkp = 10;
reg         inClk         = 1'b0;

always
begin
    #(inClkp/2) inClk = !inClk;
end

/////////////////////////////////////////

reg	[7:0] 	inRoundNumber = 8'd0;
reg	[1599:0] inData = 1600'b0;
wire	[1599:0] outData;

keccakP keccakp(.inRoundNumber(inRoundNumber), .inData(inData), .outData(outData));
 
always
begin
	inRoundNumber = 8'd0; inData = 1600'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001997b5853;
	#(inClkp);
	$stop;
end
 endmodule
